module top_module ( 
    input clk, 
    input [7:0] d, 
    input [1:0] sel, 
    output [7:0] q 
);
    wire [7:0] q1, q2, q3;
    my_dff8 inst1( .clk(clk), .d(d), .q(q1) );
    my_dff8 inst2( .clk(clk), .d(q1), .q(q2) );
    my_dff8 inst3( .clk(clk), .d(q2), .q(q3) );
    assign q = (sel == 2'b00)? d: (sel == 2'b01)? q1: (sel == 2'b10)? q2: q3;
    //always@(*) begin
//        if (sel == 00) q = d;
//    else if (sel == 01) q = q1;
//    else if (sel == 11) q = q3;
//    else q = q2;
      //  case (sel) //begin
         //   2'b00: q = d;
         //   2'b01: q = q1;
        //    2'b10: q = q2;
        //    2'b11: q = q3;
      //  endcase
    //end
endmodule
